module InstructionMemory(Address, Instruction);
	input [31:0] Address;
	output reg [31:0] Instruction;
	
	always @(*)
	begin
        //for exception test
		/*case (Address[9:2])
			8'd0:    Instruction <= 32'h08000003;
			8'd1:    Instruction <= 32'h08000008;
			8'd2:    Instruction <= 32'h08000009;
			8'd3:    Instruction <= 32'h20040003;
			8'd4:    Instruction <= 32'h20010002;
			8'd5:    Instruction <= 32'h70812002;
			8'd6:    Instruction <= 32'h20840002;
			8'd7:    Instruction <= 32'h1000ffff;
			8'd8:    Instruction <= 32'h00000000;
			8'd9:    Instruction <= 32'h20840001;
			8'd10:    Instruction <= 32'h03400008;
			default: Instruction <= 32'h0;
		endcase*/
		//for fluidity test
		/*
		case (Address[9:2])
			8'd0:    Instruction <= 32'h08000003;
			8'd1:    Instruction <= 32'h08000015;
			8'd2:    Instruction <= 32'h08000016;
			8'd3:    Instruction <= 32'h20040003;
			8'd4:    Instruction <= 32'h0c000006;
			8'd5:    Instruction <= 32'h1000ffff;
			8'd6:    Instruction <= 32'h23bdfff8;
			8'd7:    Instruction <= 32'hafbf0004;
			8'd8:    Instruction <= 32'hafa40000;
			8'd9:    Instruction <= 32'h28880001;
			8'd10:    Instruction <= 32'h11000003;
			8'd11:    Instruction <= 32'h00001026;
			8'd12:    Instruction <= 32'h23bd0008;
			8'd13:    Instruction <= 32'h03e00008;
			8'd14:    Instruction <= 32'h2084ffff;
			8'd15:    Instruction <= 32'h0c000006;
			8'd16:    Instruction <= 32'h8fa40000;
			8'd17:    Instruction <= 32'h8fbf0004;
			8'd18:   Instruction <= 32'h23bd0008;
			8'd19:   Instruction <= 32'h00821020;
			8'd20:   Instruction <= 32'h03e00008;
			8'd21:   Instruction <= 32'h1000ffff;
			8'd22:   Instruction <= 32'h1000ffff;
			default: Instruction <= 32'h0;
		endcase
		*/
		// for save-load test
		/*case (Address[9:2])
			8'd0:    Instruction <= 32'h08000003;
			8'd1:    Instruction <= 32'h0800000a;
			8'd2:    Instruction <= 32'h0800000b;
			8'd3:    Instruction <= 32'h3c083000;
			8'd4:    Instruction <= 32'h00002020;
			8'd5:    Instruction <= 32'h8d090000;
			8'd6:    Instruction <= 32'h8d0a0004;
			8'd7:    Instruction <= 32'hac890000;
			8'd8:    Instruction <= 32'hac8a0004;
			8'd9:    Instruction <= 32'h1000ffff;
			8'd10:    Instruction <= 32'h1000ffff;
			8'd11:    Instruction <= 32'h1000ffff;
			default: Instruction <= 32'h0;
		endcase*/
		//test msort
		/*case (Address[9:2])
            8'd0:Instruction <= 32'h08000003;
            8'd1:Instruction <= 32'h08000071;
            8'd2:Instruction <= 32'h08000072;
            8'd3:Instruction <= 32'h0000d820;
            8'd4:Instruction <= 32'h3c103000;
            8'd5:Instruction <= 32'h8e110000;
            8'd6:Instruction <= 32'haf600004;
            8'd7:Instruction <= 32'h001b9021;
            8'd8:Instruction <= 32'h00124821;
            8'd9:Instruction <= 32'h24080001;
            8'd10:Instruction <= 32'h237b0008;
            8'd11:Instruction <= 32'haf600004;
            8'd12:Instruction <= 32'had3b0004;
            8'd13:Instruction <= 32'h001b4821;
            8'd14:Instruction <= 32'h00085880;
            8'd15:Instruction <= 32'h01705820;
            8'd16:Instruction <= 32'h8d6a0000;
            8'd17:Instruction <= 32'had2a0000;
            8'd18:Instruction <= 32'h25080001;
            8'd19:Instruction <= 32'h0228082a;
            8'd20:Instruction <= 32'h1020fff5;
            8'd21:Instruction <= 32'h8e440004;
            8'd22:Instruction <= 32'h10800055;
            8'd23:Instruction <= 32'h0c00003e;
            8'd24:Instruction <= 32'hae420004;
            8'd25:Instruction <= 32'h0800006c;
            8'd26:Instruction <= 32'h00044821;
            8'd27:Instruction <= 32'h00055021;
            8'd28:Instruction <= 32'h237b0008;
            8'd29:Instruction <= 32'haf690004;
            8'd30:Instruction <= 32'h001b4021;
            8'd31:Instruction <= 32'h001b4821;
            8'd32:Instruction <= 32'h8d2b0000;
            8'd33:Instruction <= 32'h8d2b0004;
            8'd34:Instruction <= 32'h11600006;
            8'd35:Instruction <= 32'h8d6b0000;
            8'd36:Instruction <= 32'h8d4c0000;
            8'd37:Instruction <= 32'h018b082a;
            8'd38:Instruction <= 32'h14200005;
            8'd39:Instruction <= 32'h8d290004;
            8'd40:Instruction <= 32'h08000021;
            8'd41:Instruction <= 32'had2a0004;
            8'd42:Instruction <= 32'h8d020004;
            8'd43:Instruction <= 32'h03e00008;
            8'd44:Instruction <= 32'h000a6021;
            8'd45:Instruction <= 32'h8d8d0004;
            8'd46:Instruction <= 32'h11a00005;
            8'd47:Instruction <= 32'h8dad0000;
            8'd48:Instruction <= 32'h016d082a;
            8'd49:Instruction <= 32'h14200002;
            8'd50:Instruction <= 32'h8d8c0004;
            8'd51:Instruction <= 32'h0800002d;
            8'd52:Instruction <= 32'h8d2b0004;
            8'd53:Instruction <= 32'h8d8d0004;
            8'd54:Instruction <= 32'had8b0004;
            8'd55:Instruction <= 32'had2a0004;
            8'd56:Instruction <= 32'h000d5021;
            8'd57:Instruction <= 32'h11400002;
            8'd58:Instruction <= 32'h000b4821;
            8'd59:Instruction <= 32'h08000021;
            8'd60:Instruction <= 32'h8d020004;
            8'd61:Instruction <= 32'h03e00008;
            8'd62:Instruction <= 32'h00044021;
            8'd63:Instruction <= 32'h8d090004;
            8'd64:Instruction <= 32'h15200002;
            8'd65:Instruction <= 32'h00041021;
            8'd66:Instruction <= 32'h03e00008;
            8'd67:Instruction <= 32'h00044821;
            8'd68:Instruction <= 32'h00045021;
            8'd69:Instruction <= 32'h8d4a0004;
            8'd70:Instruction <= 32'h11400006;
            8'd71:Instruction <= 32'h8d4a0004;
            8'd72:Instruction <= 32'h11400004;
            8'd73:Instruction <= 32'h8d290004;
            8'd74:Instruction <= 32'h8d4a0004;
            8'd75:Instruction <= 32'h11400001;
            8'd76:Instruction <= 32'h08000047;
            8'd77:Instruction <= 32'h8d2a0004;
            8'd78:Instruction <= 32'had200004;
            8'd79:Instruction <= 32'h00082021;
            8'd80:Instruction <= 32'h20010008;
            8'd81:Instruction <= 32'h03a1e822;
            8'd82:Instruction <= 32'hafbf0000;
            8'd83:Instruction <= 32'hafaa0004;
            8'd84:Instruction <= 32'h0c00003e;
            8'd85:Instruction <= 32'h00025821;
            8'd86:Instruction <= 32'h8fbf0000;
            8'd87:Instruction <= 32'h8faa0004;
            8'd88:Instruction <= 32'h23bd0008;
            8'd89:Instruction <= 32'h000a2021;
            8'd90:Instruction <= 32'h20010008;
            8'd91:Instruction <= 32'h03a1e822;
            8'd92:Instruction <= 32'hafbf0000;
            8'd93:Instruction <= 32'hafab0004;
            8'd94:Instruction <= 32'h0c00003e;
            8'd95:Instruction <= 32'h00026021;
            8'd96:Instruction <= 32'h8fbf0000;
            8'd97:Instruction <= 32'h8fab0004;
            8'd98:Instruction <= 32'h23bd0008;
            8'd99:Instruction <= 32'h000b2021;
            8'd100:Instruction <= 32'h000c2821;
            8'd101:Instruction <= 32'h20010004;
            8'd102:Instruction <= 32'h03a1e822;
            8'd103:Instruction <= 32'hafbf0000;
            8'd104:Instruction <= 32'h0c00001a;
            8'd105:Instruction <= 32'h8fbf0000;
            8'd106:Instruction <= 32'h23bd0004;
            8'd107:Instruction <= 32'h03e00008;
            8'd108:Instruction <= 32'h8e480004;
            8'd109:Instruction <= 32'h8d090000;
            8'd110:Instruction <= 32'h8d080004;
            8'd111:Instruction <= 32'h1500fffd;
            8'd112:Instruction <= 32'h1000ffff;
            8'd113:Instruction <= 32'h1000ffff;
            8'd114:Instruction <= 32'h1000ffff;
            default: Instruction <= 32'h00000000;
		endcase*/
		//test interruption
		/*case(Address[9:2])
            8'd0:Instruction <= 32'h08000003;
            8'd1:Instruction <= 32'h0800002a;
            8'd2:Instruction <= 32'h08000090;
            8'd3:Instruction <= 32'h3c014000;
            8'd4:Instruction <= 32'h34210014;
            8'd5:Instruction <= 32'h00014020;
            8'd6:Instruction <= 32'h8d1c0000;
            8'd7:Instruction <= 32'h20040003;
            8'd8:Instruction <= 32'h0c00001b;
            8'd9:Instruction <= 32'h3c014000;
            8'd10:Instruction <= 32'h34210014;
            8'd11:Instruction <= 32'h00014020;
            8'd12:Instruction <= 32'h8d090000;
            8'd13:Instruction <= 32'h013ce022;
            8'd14:Instruction <= 32'h00009020;
            8'd15:Instruction <= 32'h3c01fffe;
            8'd16:Instruction <= 32'h3421c77f;
            8'd17:Instruction <= 32'h00018020;
            8'd18:Instruction <= 32'h3c014000;
            8'd19:Instruction <= 32'h34210000;
            8'd20:Instruction <= 32'h00018820;
            8'd21:Instruction <= 32'hae300000;
            8'd22:Instruction <= 32'h20100003;
            8'd23:Instruction <= 32'h20130fff;
            8'd24:Instruction <= 32'hae300008;
            8'd25:Instruction <= 32'h1000ffff;
            8'd26:Instruction <= 32'h1000ffff;
            8'd27:Instruction <= 32'h23bdfff8;
            8'd28:Instruction <= 32'hafbf0004;
            8'd29:Instruction <= 32'hafa40000;
            8'd30:Instruction <= 32'h28880001;
            8'd31:Instruction <= 32'h11000003;
            8'd32:Instruction <= 32'h00001026;
            8'd33:Instruction <= 32'h23bd0008;
            8'd34:Instruction <= 32'h03e00008;
            8'd35:Instruction <= 32'h2084ffff;
            8'd36:Instruction <= 32'h0c00001b;
            8'd37:Instruction <= 32'h8fa40000;
            8'd38:Instruction <= 32'h8fbf0004;
            8'd39:Instruction <= 32'h23bd0008;
            8'd40:Instruction <= 32'h00821020;
            8'd41:Instruction <= 32'h03e00008;
            8'd42:Instruction <= 32'h32100000;
            8'd43:Instruction <= 32'hae300008;
            8'd44:Instruction <= 32'h200107d0;
            8'd45:Instruction <= 32'h0032082a;
            8'd46:Instruction <= 32'h1420005f;
            8'd47:Instruction <= 32'h32690f00;
            8'd48:Instruction <= 32'h36730f00;
            8'd49:Instruction <= 32'h20010e00;
            8'd50:Instruction <= 32'h10290007;
            8'd51:Instruction <= 32'h20010d00;
            8'd52:Instruction <= 32'h10290008;
            8'd53:Instruction <= 32'h20010b00;
            8'd54:Instruction <= 32'h10290009;
            8'd55:Instruction <= 32'h20010700;
            8'd56:Instruction <= 32'h1029000a;
            8'd57:Instruction <= 32'h08000043;
            8'd58:Instruction <= 32'h32730dff;
            8'd59:Instruction <= 32'h001c2102;
            8'd60:Instruction <= 32'h08000046;
            8'd61:Instruction <= 32'h32730bff;
            8'd62:Instruction <= 32'h001c2202;
            8'd63:Instruction <= 32'h08000046;
            8'd64:Instruction <= 32'h327307ff;
            8'd65:Instruction <= 32'h001c2302;
            8'd66:Instruction <= 32'h08000046;
            8'd67:Instruction <= 32'h32730eff;
            8'd68:Instruction <= 32'h001c2002;
            8'd69:Instruction <= 32'h08000046;
            8'd70:Instruction <= 32'h367300ff;
            8'd71:Instruction <= 32'h3084000f;
            8'd72:Instruction <= 32'h20010000;
            8'd73:Instruction <= 32'h1024001f;
            8'd74:Instruction <= 32'h20010001;
            8'd75:Instruction <= 32'h1024001f;
            8'd76:Instruction <= 32'h20010002;
            8'd77:Instruction <= 32'h1024001f;
            8'd78:Instruction <= 32'h20010003;
            8'd79:Instruction <= 32'h1024001f;
            8'd80:Instruction <= 32'h20010004;
            8'd81:Instruction <= 32'h1024001f;
            8'd82:Instruction <= 32'h20010005;
            8'd83:Instruction <= 32'h1024001f;
            8'd84:Instruction <= 32'h20010006;
            8'd85:Instruction <= 32'h1024001f;
            8'd86:Instruction <= 32'h20010007;
            8'd87:Instruction <= 32'h1024001f;
            8'd88:Instruction <= 32'h20010008;
            8'd89:Instruction <= 32'h1024001f;
            8'd90:Instruction <= 32'h20010009;
            8'd91:Instruction <= 32'h1024001f;
            8'd92:Instruction <= 32'h2001000a;
            8'd93:Instruction <= 32'h1024001f;
            8'd94:Instruction <= 32'h2001000b;
            8'd95:Instruction <= 32'h1024001f;
            8'd96:Instruction <= 32'h2001000c;
            8'd97:Instruction <= 32'h1024001f;
            8'd98:Instruction <= 32'h2001000d;
            8'd99:Instruction <= 32'h1024001f;
            8'd100:Instruction <= 32'h2001000e;
            8'd101:Instruction <= 32'h1024001f;
            8'd102:Instruction <= 32'h2001000f;
            8'd103:Instruction <= 32'h1024001f;
            8'd104:Instruction <= 32'h08000089;
            8'd105:Instruction <= 32'h32730f40;
            8'd106:Instruction <= 32'h08000089;
            8'd107:Instruction <= 32'h32730f79;
            8'd108:Instruction <= 32'h08000089;
            8'd109:Instruction <= 32'h32730f24;
            8'd110:Instruction <= 32'h08000089;
            8'd111:Instruction <= 32'h32730f30;
            8'd112:Instruction <= 32'h08000089;
            8'd113:Instruction <= 32'h32730f19;
            8'd114:Instruction <= 32'h08000089;
            8'd115:Instruction <= 32'h32730f12;
            8'd116:Instruction <= 32'h08000089;
            8'd117:Instruction <= 32'h32730f02;
            8'd118:Instruction <= 32'h08000089;
            8'd119:Instruction <= 32'h32730f78;
            8'd120:Instruction <= 32'h08000089;
            8'd121:Instruction <= 32'h32730f00;
            8'd122:Instruction <= 32'h08000089;
            8'd123:Instruction <= 32'h32730f10;
            8'd124:Instruction <= 32'h08000089;
            8'd125:Instruction <= 32'h32730f08;
            8'd126:Instruction <= 32'h08000089;
            8'd127:Instruction <= 32'h32730f03;
            8'd128:Instruction <= 32'h08000089;
            8'd129:Instruction <= 32'h32730f46;
            8'd130:Instruction <= 32'h08000089;
            8'd131:Instruction <= 32'h32730f21;
            8'd132:Instruction <= 32'h08000089;
            8'd133:Instruction <= 32'h32730f06;
            8'd134:Instruction <= 32'h08000089;
            8'd135:Instruction <= 32'h32730f0e;
            8'd136:Instruction <= 32'h08000089;
            8'd137:Instruction <= 32'hae330010;
            8'd138:Instruction <= 32'h22520001;
            8'd139:Instruction <= 32'h36100003;
            8'd140:Instruction <= 32'hae300008;
            8'd141:Instruction <= 32'h03400008;
            8'd142:Instruction <= 32'h0002e020;
            8'd143:Instruction <= 32'h0800002f;
            8'd144:Instruction <= 32'h1000ffff;
            default: Instruction<=32'h0;
		endcase*/
		//MSORT FINAL
		case(Address[9:2])
			8'd0:Instruction <= 32'h08000003;
			8'd1:Instruction <= 32'h08000082;
			8'd2:Instruction <= 32'h080000ea;
			8'd3:Instruction <= 32'h3c014000;
			8'd4:Instruction <= 32'h34210014;
			8'd5:Instruction <= 32'h00014020;
			8'd6:Instruction <= 32'h8d1c0000;
			8'd7:Instruction <= 32'h0000d820;
			8'd8:Instruction <= 32'h3c103000;
			8'd9:Instruction <= 32'h8e110000;
			8'd10:Instruction <= 32'haf600004;
			8'd11:Instruction <= 32'h001b9021;
			8'd12:Instruction <= 32'h00124821;
			8'd13:Instruction <= 32'h24080001;
			8'd14:Instruction <= 32'h237b0008;
			8'd15:Instruction <= 32'haf600004;
			8'd16:Instruction <= 32'had3b0004;
			8'd17:Instruction <= 32'h001b4821;
			8'd18:Instruction <= 32'h00085880;
			8'd19:Instruction <= 32'h01705820;
			8'd20:Instruction <= 32'h8d6a0000;
			8'd21:Instruction <= 32'had2a0000;
			8'd22:Instruction <= 32'h25080001;
			8'd23:Instruction <= 32'h0228082a;
			8'd24:Instruction <= 32'h1020fff5;
			8'd25:Instruction <= 32'h8e440004;
			8'd26:Instruction <= 32'h10800055;
			8'd27:Instruction <= 32'h0c000042;
			8'd28:Instruction <= 32'hae420004;
			8'd29:Instruction <= 32'h08000070;
			8'd30:Instruction <= 32'h00044821;
			8'd31:Instruction <= 32'h00055021;
			8'd32:Instruction <= 32'h237b0008;
			8'd33:Instruction <= 32'haf690004;
			8'd34:Instruction <= 32'h001b4021;
			8'd35:Instruction <= 32'h001b4821;
			8'd36:Instruction <= 32'h8d2b0000;
			8'd37:Instruction <= 32'h8d2b0004;
			8'd38:Instruction <= 32'h11600006;
			8'd39:Instruction <= 32'h8d6b0000;
			8'd40:Instruction <= 32'h8d4c0000;
			8'd41:Instruction <= 32'h018b082a;
			8'd42:Instruction <= 32'h14200005;
			8'd43:Instruction <= 32'h8d290004;
			8'd44:Instruction <= 32'h08000025;
			8'd45:Instruction <= 32'had2a0004;
			8'd46:Instruction <= 32'h8d020004;
			8'd47:Instruction <= 32'h03e00008;
			8'd48:Instruction <= 32'h000a6021;
			8'd49:Instruction <= 32'h8d8d0004;
			8'd50:Instruction <= 32'h11a00005;
			8'd51:Instruction <= 32'h8dad0000;
			8'd52:Instruction <= 32'h016d082a;
			8'd53:Instruction <= 32'h14200002;
			8'd54:Instruction <= 32'h8d8c0004;
			8'd55:Instruction <= 32'h08000031;
			8'd56:Instruction <= 32'h8d2b0004;
			8'd57:Instruction <= 32'h8d8d0004;
			8'd58:Instruction <= 32'had8b0004;
			8'd59:Instruction <= 32'had2a0004;
			8'd60:Instruction <= 32'h000d5021;
			8'd61:Instruction <= 32'h11400002;
			8'd62:Instruction <= 32'h000b4821;
			8'd63:Instruction <= 32'h08000025;
			8'd64:Instruction <= 32'h8d020004;
			8'd65:Instruction <= 32'h03e00008;
			8'd66:Instruction <= 32'h00044021;
			8'd67:Instruction <= 32'h8d090004;
			8'd68:Instruction <= 32'h15200002;
			8'd69:Instruction <= 32'h00041021;
			8'd70:Instruction <= 32'h03e00008;
			8'd71:Instruction <= 32'h00044821;
			8'd72:Instruction <= 32'h00045021;
			8'd73:Instruction <= 32'h8d4a0004;
			8'd74:Instruction <= 32'h11400006;
			8'd75:Instruction <= 32'h8d4a0004;
			8'd76:Instruction <= 32'h11400004;
			8'd77:Instruction <= 32'h8d290004;
			8'd78:Instruction <= 32'h8d4a0004;
			8'd79:Instruction <= 32'h11400001;
			8'd80:Instruction <= 32'h0800004b;
			8'd81:Instruction <= 32'h8d2a0004;
			8'd82:Instruction <= 32'had200004;
			8'd83:Instruction <= 32'h00082021;
			8'd84:Instruction <= 32'h20010008;
			8'd85:Instruction <= 32'h03a1e822;
			8'd86:Instruction <= 32'hafbf0000;
			8'd87:Instruction <= 32'hafaa0004;
			8'd88:Instruction <= 32'h0c000042;
			8'd89:Instruction <= 32'h00025821;
			8'd90:Instruction <= 32'h8fbf0000;
			8'd91:Instruction <= 32'h8faa0004;
			8'd92:Instruction <= 32'h23bd0008;
			8'd93:Instruction <= 32'h000a2021;
			8'd94:Instruction <= 32'h20010008;
			8'd95:Instruction <= 32'h03a1e822;
			8'd96:Instruction <= 32'hafbf0000;
			8'd97:Instruction <= 32'hafab0004;
			8'd98:Instruction <= 32'h0c000042;
			8'd99:Instruction <= 32'h00026021;
			8'd100:Instruction <= 32'h8fbf0000;
			8'd101:Instruction <= 32'h8fab0004;
			8'd102:Instruction <= 32'h23bd0008;
			8'd103:Instruction <= 32'h000b2021;
			8'd104:Instruction <= 32'h000c2821;
			8'd105:Instruction <= 32'h20010004;
			8'd106:Instruction <= 32'h03a1e822;
			8'd107:Instruction <= 32'hafbf0000;
			8'd108:Instruction <= 32'h0c00001e;
			8'd109:Instruction <= 32'h8fbf0000;
			8'd110:Instruction <= 32'h23bd0004;
			8'd111:Instruction <= 32'h03e00008;
			8'd112:Instruction <= 32'h8c180000;
			8'd113:Instruction <= 32'h3c014000;
			8'd114:Instruction <= 32'h34210014;
			8'd115:Instruction <= 32'h00014020;
			8'd116:Instruction <= 32'h8d090000;
			8'd117:Instruction <= 32'h013ce022;
			8'd118:Instruction <= 32'h00009020;
			8'd119:Instruction <= 32'h3c01fffe;
			8'd120:Instruction <= 32'h3421c77f;
			8'd121:Instruction <= 32'h00018020;
			8'd122:Instruction <= 32'h3c014000;
			8'd123:Instruction <= 32'h34210000;
			8'd124:Instruction <= 32'h00018820;
			8'd125:Instruction <= 32'hae300000;
			8'd126:Instruction <= 32'h20100003;
			8'd127:Instruction <= 32'h20130fff;
			8'd128:Instruction <= 32'hae300008;
			8'd129:Instruction <= 32'h1000ffff;
			8'd130:Instruction <= 32'h32100000;
			8'd131:Instruction <= 32'hae300008;
			8'd132:Instruction <= 32'h200107d0;
			8'd133:Instruction <= 32'h0032082a;
			8'd134:Instruction <= 32'h1420005f;
			8'd135:Instruction <= 32'h32690f00;
			8'd136:Instruction <= 32'h36730f00;
			8'd137:Instruction <= 32'h20010e00;
			8'd138:Instruction <= 32'h10290007;
			8'd139:Instruction <= 32'h20010d00;
			8'd140:Instruction <= 32'h10290008;
			8'd141:Instruction <= 32'h20010b00;
			8'd142:Instruction <= 32'h10290009;
			8'd143:Instruction <= 32'h20010700;
			8'd144:Instruction <= 32'h1029000a;
			8'd145:Instruction <= 32'h0800009b;
			8'd146:Instruction <= 32'h32730dff;
			8'd147:Instruction <= 32'h001c2102;
			8'd148:Instruction <= 32'h0800009e;
			8'd149:Instruction <= 32'h32730bff;
			8'd150:Instruction <= 32'h001c2202;
			8'd151:Instruction <= 32'h0800009e;
			8'd152:Instruction <= 32'h327307ff;
			8'd153:Instruction <= 32'h001c2302;
			8'd154:Instruction <= 32'h0800009e;
			8'd155:Instruction <= 32'h32730eff;
			8'd156:Instruction <= 32'h001c2002;
			8'd157:Instruction <= 32'h0800009e;
			8'd158:Instruction <= 32'h367300ff;
			8'd159:Instruction <= 32'h3084000f;
			8'd160:Instruction <= 32'h20010000;
			8'd161:Instruction <= 32'h1024001f;
			8'd162:Instruction <= 32'h20010001;
			8'd163:Instruction <= 32'h1024001f;
			8'd164:Instruction <= 32'h20010002;
			8'd165:Instruction <= 32'h1024001f;
			8'd166:Instruction <= 32'h20010003;
			8'd167:Instruction <= 32'h1024001f;
			8'd168:Instruction <= 32'h20010004;
			8'd169:Instruction <= 32'h1024001f;
			8'd170:Instruction <= 32'h20010005;
			8'd171:Instruction <= 32'h1024001f;
			8'd172:Instruction <= 32'h20010006;
			8'd173:Instruction <= 32'h1024001f;
			8'd174:Instruction <= 32'h20010007;
			8'd175:Instruction <= 32'h1024001f;
			8'd176:Instruction <= 32'h20010008;
			8'd177:Instruction <= 32'h1024001f;
			8'd178:Instruction <= 32'h20010009;
			8'd179:Instruction <= 32'h1024001f;
			8'd180:Instruction <= 32'h2001000a;
			8'd181:Instruction <= 32'h1024001f;
			8'd182:Instruction <= 32'h2001000b;
			8'd183:Instruction <= 32'h1024001f;
			8'd184:Instruction <= 32'h2001000c;
			8'd185:Instruction <= 32'h1024001f;
			8'd186:Instruction <= 32'h2001000d;
			8'd187:Instruction <= 32'h1024001f;
			8'd188:Instruction <= 32'h2001000e;
			8'd189:Instruction <= 32'h1024001f;
			8'd190:Instruction <= 32'h2001000f;
			8'd191:Instruction <= 32'h1024001f;
			8'd192:Instruction <= 32'h080000e1;
			8'd193:Instruction <= 32'h32730f40;
			8'd194:Instruction <= 32'h080000e1;
			8'd195:Instruction <= 32'h32730f79;
			8'd196:Instruction <= 32'h080000e1;
			8'd197:Instruction <= 32'h32730f24;
			8'd198:Instruction <= 32'h080000e1;
			8'd199:Instruction <= 32'h32730f30;
			8'd200:Instruction <= 32'h080000e1;
			8'd201:Instruction <= 32'h32730f19;
			8'd202:Instruction <= 32'h080000e1;
			8'd203:Instruction <= 32'h32730f12;
			8'd204:Instruction <= 32'h080000e1;
			8'd205:Instruction <= 32'h32730f02;
			8'd206:Instruction <= 32'h080000e1;
			8'd207:Instruction <= 32'h32730f78;
			8'd208:Instruction <= 32'h080000e1;
			8'd209:Instruction <= 32'h32730f00;
			8'd210:Instruction <= 32'h080000e1;
			8'd211:Instruction <= 32'h32730f10;
			8'd212:Instruction <= 32'h080000e1;
			8'd213:Instruction <= 32'h32730f08;
			8'd214:Instruction <= 32'h080000e1;
			8'd215:Instruction <= 32'h32730f03;
			8'd216:Instruction <= 32'h080000e1;
			8'd217:Instruction <= 32'h32730f46;
			8'd218:Instruction <= 32'h080000e1;
			8'd219:Instruction <= 32'h32730f21;
			8'd220:Instruction <= 32'h080000e1;
			8'd221:Instruction <= 32'h32730f06;
			8'd222:Instruction <= 32'h080000e1;
			8'd223:Instruction <= 32'h32730f0e;
			8'd224:Instruction <= 32'h080000e1;
			8'd225:Instruction <= 32'hae330010;
			8'd226:Instruction <= 32'h22520001;
			8'd227:Instruction <= 32'h36100003;
			8'd228:Instruction <= 32'hae300008;
			8'd229:Instruction <= 32'h03400008;
			8'd230:Instruction <= 32'h8f1c0000;
			8'd231:Instruction <= 32'h00009020;
			8'd232:Instruction <= 32'h8f180004;
			8'd233:Instruction <= 32'h08000087;
			8'd234:Instruction <= 32'h1000ffff;
			default: Instruction<=32'h0;
		endcase
	end	
endmodule
